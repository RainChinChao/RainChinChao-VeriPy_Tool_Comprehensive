module else_self_gen_290( input clk, input reset, input [31:0]array_ref_m_wire_0, output [31:0]segment_0); 
	wire [31:0]segment_0;
	//Proceed with segment_0 = array_ref_m_wire_0
	delay Value_HDL_0 ( clk, reset, array_ref_m_wire_0, segment_0);
endmodule