module If__V_1_if_calculation(input [31:0]input_bit, input [31:0]zero, input [31:0]array_ref_wire_1, input [31:0]array_ref_m_wire_1, output [31:0]segment_1, input clk, input reset);



	//Proceed with segment_1 = delay(array_ref_wire_1) 
	wire [31:0]segment_1;
	delay Value_HDL_Level0_1 ( clk, reset, array_ref_wire_1, segment_1);




endmodule
