module else_self_gen_279( input clk, input reset, input [31:0]array_ref_m_wire_9, output [31:0]segment_9); 
	wire [31:0]segment_9;
	//Proceed with segment_9 = array_ref_m_wire_9
	delay Value_HDL_0 ( clk, reset, array_ref_m_wire_9, segment_9);
endmodule