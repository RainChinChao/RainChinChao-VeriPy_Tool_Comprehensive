`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.12.2024 13:36:34
// Design Name: 
// Module Name: toptop
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




//module toptop( input [31:0]a, input [31:0]b, output [31:0]temp_real_31, output [31:0]temp_imag_31, input clk

//    );
    
    
//reg [31:0]X_real_0;
//reg [31:0]X_imag_0;
//always @(posedge clk) begin 
//	X_real_0 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_0 <= a;
//end
//reg [31:0]X_real_1;
//reg [31:0]X_imag_1;
//always @(posedge clk) begin 
//	X_real_1 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_1 <= a;
//end
//reg [31:0]X_real_2;
//reg [31:0]X_imag_2;
//always @(posedge clk) begin 
//	X_real_2 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_2 <= a;
//end
//reg [31:0]X_real_3;
//reg [31:0]X_imag_3;
//always @(posedge clk) begin 
//	X_real_3 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_3 <= a;
//end
//reg [31:0]X_real_4;
//reg [31:0]X_imag_4;
//always @(posedge clk) begin 
//	X_real_4 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_4 <= a;
//end
//reg [31:0]X_real_5;
//reg [31:0]X_imag_5;
//always @(posedge clk) begin 
//	X_real_5 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_5 <= a;
//end
//reg [31:0]X_real_6;
//reg [31:0]X_imag_6;
//always @(posedge clk) begin 
//	X_real_6 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_6 <= a;
//end
//reg [31:0]X_real_7;
//reg [31:0]X_imag_7;
//always @(posedge clk) begin 
//	X_real_7 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_7 <= a;
//end
//reg [31:0]X_real_8;
//reg [31:0]X_imag_8;
//always @(posedge clk) begin 
//	X_real_8 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_8 <= a;
//end
//reg [31:0]X_real_9;
//reg [31:0]X_imag_9;
//always @(posedge clk) begin 
//	X_real_9 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_9 <= a;
//end
//reg [31:0]X_real_10;
//reg [31:0]X_imag_10;
//always @(posedge clk) begin 
//	X_real_10 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_10 <= a;
//end
//reg [31:0]X_real_11;
//reg [31:0]X_imag_11;
//always @(posedge clk) begin 
//	X_real_11 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_11 <= a;
//end
//reg [31:0]X_real_12;
//reg [31:0]X_imag_12;
//always @(posedge clk) begin 
//	X_real_12 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_12 <= a;
//end
//reg [31:0]X_real_13;
//reg [31:0]X_imag_13;
//always @(posedge clk) begin 
//	X_real_13 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_13 <= a;
//end
//reg [31:0]X_real_14;
//reg [31:0]X_imag_14;
//always @(posedge clk) begin 
//	X_real_14 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_14 <= a;
//end
//reg [31:0]X_real_15;
//reg [31:0]X_imag_15;
//always @(posedge clk) begin 
//	X_real_15 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_15 <= a;
//end
//reg [31:0]X_real_16;
//reg [31:0]X_imag_16;
//always @(posedge clk) begin 
//	X_real_16 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_16 <= a;
//end
//reg [31:0]X_real_17;
//reg [31:0]X_imag_17;
//always @(posedge clk) begin 
//	X_real_17 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_17 <= a;
//end
//reg [31:0]X_real_18;
//reg [31:0]X_imag_18;
//always @(posedge clk) begin 
//	X_real_18 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_18 <= a;
//end
//reg [31:0]X_real_19;
//reg [31:0]X_imag_19;
//always @(posedge clk) begin 
//	X_real_19 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_19 <= a;
//end
//reg [31:0]X_real_20;
//reg [31:0]X_imag_20;
//always @(posedge clk) begin 
//	X_real_20 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_20 <= a;
//end
//reg [31:0]X_real_21;
//reg [31:0]X_imag_21;
//always @(posedge clk) begin 
//	X_real_21 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_21 <= a;
//end
//reg [31:0]X_real_22;
//reg [31:0]X_imag_22;
//always @(posedge clk) begin 
//	X_real_22 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_22 <= a;
//end
//reg [31:0]X_real_23;
//reg [31:0]X_imag_23;
//always @(posedge clk) begin 
//	X_real_23 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_23 <= a;
//end
//reg [31:0]X_real_24;
//reg [31:0]X_imag_24;
//always @(posedge clk) begin 
//	X_real_24 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_24 <= a;
//end
//reg [31:0]X_real_25;
//reg [31:0]X_imag_25;
//always @(posedge clk) begin 
//	X_real_25 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_25 <= a;
//end
//reg [31:0]X_real_26;
//reg [31:0]X_imag_26;
//always @(posedge clk) begin 
//	X_real_26 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_26 <= a;
//end
//reg [31:0]X_real_27;
//reg [31:0]X_imag_27;
//always @(posedge clk) begin 
//	X_real_27 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_27 <= a;
//end
//reg [31:0]X_real_28;
//reg [31:0]X_imag_28;
//always @(posedge clk) begin 
//	X_real_28 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_28 <= a;
//end
//reg [31:0]X_real_29;
//reg [31:0]X_imag_29;
//always @(posedge clk) begin 
//	X_real_29 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_29 <= a;
//end
//reg [31:0]X_real_30;
//reg [31:0]X_imag_30;
//always @(posedge clk) begin 
//	X_real_30 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_30 <= a;
//end
//reg [31:0]X_real_31;
//reg [31:0]X_imag_31;
//always @(posedge clk) begin 
//	X_real_31 <= a;
//end
//always @(posedge clk) begin 
//	X_imag_31 <= a;
//end
    
//    top tt2( X_real_0, X_imag_0, X_real_1, X_imag_1, X_real_2, X_imag_2, X_real_3, X_imag_3, X_real_4, X_imag_4, X_real_5, X_imag_5, X_real_6, X_imag_6, X_real_7, X_imag_7, X_real_8, X_imag_8, X_real_9, X_imag_9, X_real_10, X_imag_10, X_real_11, X_imag_11, X_real_12, X_imag_12, X_real_13, X_imag_13, X_real_14, X_imag_14, X_real_15, X_imag_15, X_real_16, X_imag_16, X_real_17, X_imag_17, X_real_18, X_imag_18, X_real_19, X_imag_19, X_real_20, X_imag_20, X_real_21, X_imag_21, X_real_22, X_imag_22, X_real_23, X_imag_23, X_real_24, X_imag_24, X_real_25, X_imag_25, X_real_26, X_imag_26, X_real_27, X_imag_27, X_real_28, X_imag_28, X_real_29, X_imag_29, X_real_30, X_imag_30, X_real_31, X_imag_31, temp_real_31,temp_imag_31, clk, start, valid, busy, reset); 

    
    
    
//endmodule
















module toptop( input [31:0]I, output [31:0]x_15,  input clk, input reset

    );

reg [31:0]X_real_0 = 0;

always @(posedge clk) begin 
	X_real_0 <= I;
end

reg [31:0]X_real_1 = 0;

always @(posedge clk) begin 
	X_real_1 <= X_real_0;
end

reg [31:0]X_real_2 = 0;

always @(posedge clk) begin 
	X_real_2 <= X_real_1;
end

reg [31:0]X_real_3 = 0;

always @(posedge clk) begin 
	X_real_3 <= X_real_2;
end

reg [31:0]X_real_4 = 0;

always @(posedge clk) begin 
	X_real_4 <= X_real_3;
end

reg [31:0]X_real_5 = 0;

always @(posedge clk) begin 
	X_real_5 <= X_real_4;
end

reg [31:0]X_real_6 = 0;

always @(posedge clk) begin 
	X_real_6 <= X_real_5;
end

reg [31:0]X_real_7 = 0;

always @(posedge clk) begin 
	X_real_7 <= X_real_6;
end

reg [31:0]X_real_8 = 0;

always @(posedge clk) begin 
	X_real_8 <= X_real_7;
end

reg [31:0]X_real_9 = 0;

always @(posedge clk) begin 
	X_real_9 <= X_real_8;
end

reg [31:0]X_real_10 = 0;

always @(posedge clk) begin 
	X_real_10 <= X_real_9;
end

reg [31:0]X_real_11 = 0;

always @(posedge clk) begin 
	X_real_11 <= X_real_10;
end

reg [31:0]X_real_12 = 0;

always @(posedge clk) begin 
	X_real_12 <= X_real_11;
end

reg [31:0]X_real_13 = 0;

always @(posedge clk) begin 
	X_real_13 <= X_real_12;
end

reg [31:0]X_real_14 = 0;

always @(posedge clk) begin 
	X_real_14 <= X_real_13;
end

reg [31:0]X_real_15 = 0;

always @(posedge clk) begin 
	X_real_15 <= X_real_14;
end






    top tt2( X_real_0, X_real_1, X_real_2, X_real_3, X_real_4, X_real_5, X_real_6, X_real_7, X_real_8, X_real_9, X_real_10, X_real_11, X_real_12, X_real_13, X_real_14, X_real_15,x_15, clk, reset); 

    
    
    
endmodule









