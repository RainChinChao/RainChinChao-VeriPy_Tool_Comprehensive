module if_self_gen_297( input clk, input reset, input [31:0]array_ref_wire_7, output [31:0]segment_7); 
	wire [31:0]segment_7;
	//Proceed with segment_7 = array_ref_wire_7
	delay Value_HDL_0 ( clk, reset, array_ref_wire_7, segment_7);
endmodule