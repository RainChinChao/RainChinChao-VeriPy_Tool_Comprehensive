module if_self_gen_293( input clk, input reset, input [31:0]array_ref_wire_3, output [31:0]segment_3); 
	wire [31:0]segment_3;
	//Proceed with segment_3 = array_ref_wire_3
	delay Value_HDL_0 ( clk, reset, array_ref_wire_3, segment_3);
endmodule