module if_self_gen_291( input clk, input reset, input [31:0]array_ref_wire_1, output [31:0]segment_1); 
	wire [31:0]segment_1;
	//Proceed with segment_1 = array_ref_wire_1
	delay Value_HDL_0 ( clk, reset, array_ref_wire_1, segment_1);
endmodule