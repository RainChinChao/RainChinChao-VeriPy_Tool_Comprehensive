module else_self_gen_298( input clk, input reset, input [31:0]array_ref_m_wire_8, output [31:0]segment_8); 
	wire [31:0]segment_8;
	//Proceed with segment_8 = array_ref_m_wire_8
	delay Value_HDL_0 ( clk, reset, array_ref_m_wire_8, segment_8);
endmodule