module if_self_gen_296( input clk, input reset, input [31:0]array_ref_wire_6, output [31:0]segment_6); 
	wire [31:0]segment_6;
	//Proceed with segment_6 = array_ref_wire_6
	delay Value_HDL_0 ( clk, reset, array_ref_wire_6, segment_6);
endmodule