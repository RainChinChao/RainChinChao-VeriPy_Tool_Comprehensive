module else_self_gen_272( input clk, input reset, input [31:0]array_ref_m_wire_2, output [31:0]segment_2); 
	wire [31:0]segment_2;
	//Proceed with segment_2 = array_ref_m_wire_2
	delay Value_HDL_0 ( clk, reset, array_ref_m_wire_2, segment_2);
endmodule