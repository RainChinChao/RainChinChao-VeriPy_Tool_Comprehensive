module If__V_9_else_calculation(input [31:0]input_bit, input [31:0]zero, input [31:0]array_ref_wire_9, input [31:0]array_ref_m_wire_9, output [31:0]segment_9, input clk, input reset, input start, output valid, output busy);



	//Proceed with segment_9 = delay(array_ref_m_wire_9) 
	wire [31:0]segment_9;
	delay Value_HDL_Level0_9 ( clk, reset, array_ref_m_wire_9, segment_9);




endmodule
