module If_test( input [31:0]input_bit, output [31:0]segment_0, output [31:0]segment_1, output [31:0]segment_2, output [31:0]segment_3, output [31:0]segment_4, output [31:0]segment_5, output [31:0]segment_6, output [31:0]segment_7, output [31:0]segment_8, output [31:0]segment_9, input clk, input reset); 



	// Generate the array ref[10]
	reg [31:0] array_ref_0 = 65536; 
	wire [31:0] array_ref_wire_0;
	assign  array_ref_wire_0 = array_ref_0;
	reg [31:0] array_ref_1 = 4294901760; 
	wire [31:0] array_ref_wire_1;
	assign  array_ref_wire_1 = array_ref_1;
	reg [31:0] array_ref_2 = 65536; 
	wire [31:0] array_ref_wire_2;
	assign  array_ref_wire_2 = array_ref_2;
	reg [31:0] array_ref_3 = 4294901760; 
	wire [31:0] array_ref_wire_3;
	assign  array_ref_wire_3 = array_ref_3;
	reg [31:0] array_ref_4 = 65536; 
	wire [31:0] array_ref_wire_4;
	assign  array_ref_wire_4 = array_ref_4;
	reg [31:0] array_ref_5 = 4294901760; 
	wire [31:0] array_ref_wire_5;
	assign  array_ref_wire_5 = array_ref_5;
	reg [31:0] array_ref_6 = 65536; 
	wire [31:0] array_ref_wire_6;
	assign  array_ref_wire_6 = array_ref_6;
	reg [31:0] array_ref_7 = 4294901760; 
	wire [31:0] array_ref_wire_7;
	assign  array_ref_wire_7 = array_ref_7;
	reg [31:0] array_ref_8 = 65536; 
	wire [31:0] array_ref_wire_8;
	assign  array_ref_wire_8 = array_ref_8;
	reg [31:0] array_ref_9 = 4294901760; 
	wire [31:0] array_ref_wire_9;
	assign  array_ref_wire_9 = array_ref_9;
	// End the array ref[10]






	// Generate the array ref_m[10]
	reg [31:0] array_ref_m_0 = 4294901760; 
	wire [31:0] array_ref_m_wire_0;
	assign  array_ref_m_wire_0 = array_ref_m_0;
	reg [31:0] array_ref_m_1 = 65536; 
	wire [31:0] array_ref_m_wire_1;
	assign  array_ref_m_wire_1 = array_ref_m_1;
	reg [31:0] array_ref_m_2 = 4294901760; 
	wire [31:0] array_ref_m_wire_2;
	assign  array_ref_m_wire_2 = array_ref_m_2;
	reg [31:0] array_ref_m_3 = 65536; 
	wire [31:0] array_ref_m_wire_3;
	assign  array_ref_m_wire_3 = array_ref_m_3;
	reg [31:0] array_ref_m_4 = 4294901760; 
	wire [31:0] array_ref_m_wire_4;
	assign  array_ref_m_wire_4 = array_ref_m_4;
	reg [31:0] array_ref_m_5 = 65536; 
	wire [31:0] array_ref_m_wire_5;
	assign  array_ref_m_wire_5 = array_ref_m_5;
	reg [31:0] array_ref_m_6 = 4294901760; 
	wire [31:0] array_ref_m_wire_6;
	assign  array_ref_m_wire_6 = array_ref_m_6;
	reg [31:0] array_ref_m_7 = 65536; 
	wire [31:0] array_ref_m_wire_7;
	assign  array_ref_m_wire_7 = array_ref_m_7;
	reg [31:0] array_ref_m_8 = 4294901760; 
	wire [31:0] array_ref_m_wire_8;
	assign  array_ref_m_wire_8 = array_ref_m_8;
	reg [31:0] array_ref_m_9 = 65536; 
	wire [31:0] array_ref_m_wire_9;
	assign  array_ref_m_wire_9 = array_ref_m_9;
	// End the array ref_m[10]




	wire [31:0]segment_0;
	//Proceed with one function if calculation.
	if_else_self_gen_290 else_HDL_290( clk , reset, input_bit, array_ref_wire_0, array_ref_m_wire_0, segment_0);





	wire [31:0]segment_1;
	//Proceed with one function if calculation.
	if_else_self_gen_291 else_HDL_291( clk , reset, input_bit, array_ref_m_wire_1, array_ref_wire_1, segment_1);





	wire [31:0]segment_2;
	//Proceed with one function if calculation.
	if_else_self_gen_292 else_HDL_292( clk , reset, input_bit, array_ref_m_wire_2, array_ref_wire_2, segment_2);





	wire [31:0]segment_3;
	//Proceed with one function if calculation.
	if_else_self_gen_293 else_HDL_293( clk , reset, input_bit, array_ref_wire_3, array_ref_m_wire_3, segment_3);





	wire [31:0]segment_4;
	//Proceed with one function if calculation.
	if_else_self_gen_294 else_HDL_294( clk , reset, input_bit, array_ref_wire_4, array_ref_m_wire_4, segment_4);





	wire [31:0]segment_5;
	//Proceed with one function if calculation.
	if_else_self_gen_295 else_HDL_295( clk , reset, input_bit, array_ref_m_wire_5, array_ref_wire_5, segment_5);





	wire [31:0]segment_6;
	//Proceed with one function if calculation.
	if_else_self_gen_296 else_HDL_296( clk , reset, input_bit, array_ref_wire_6, array_ref_m_wire_6, segment_6);





	wire [31:0]segment_7;
	//Proceed with one function if calculation.
	if_else_self_gen_297 else_HDL_297( clk , reset, input_bit, array_ref_wire_7, array_ref_m_wire_7, segment_7);





	wire [31:0]segment_8;
	//Proceed with one function if calculation.
	if_else_self_gen_298 else_HDL_298( clk , reset, input_bit, array_ref_wire_8, array_ref_m_wire_8, segment_8);





	wire [31:0]segment_9;
	//Proceed with one function if calculation.
	if_else_self_gen_299 else_HDL_299( clk , reset, input_bit, array_ref_wire_9, array_ref_m_wire_9, segment_9);





endmodule