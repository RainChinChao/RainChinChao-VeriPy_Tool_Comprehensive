module if_self_gen_294( input clk, input reset, input [31:0]array_ref_wire_4, output [31:0]segment_4); 
	wire [31:0]segment_4;
	//Proceed with segment_4 = array_ref_wire_4
	delay Value_HDL_0 ( clk, reset, array_ref_wire_4, segment_4);
endmodule