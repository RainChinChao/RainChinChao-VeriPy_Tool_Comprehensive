module If__V_6_if_calculation(input [31:0]input_bit, input [31:0]zero, input [31:0]array_ref_wire_6, input [31:0]array_ref_m_wire_6, output [31:0]segment_6, input clk, input reset);



	//Proceed with segment_6 = delay(array_ref_wire_6) 
	wire [31:0]segment_6;
	delay Value_HDL_Level0_6 ( clk, reset, array_ref_wire_6, segment_6);




endmodule
