module if_self_gen_295( input clk, input reset, input [31:0]array_ref_wire_5, output [31:0]segment_5); 
	wire [31:0]segment_5;
	//Proceed with segment_5 = array_ref_wire_5
	delay Value_HDL_0 ( clk, reset, array_ref_wire_5, segment_5);
endmodule